* /home/edeelep/eSim-Workspace/sc_test/sc_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu 10 Mar 2022 09:52:14 AM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  clk Net-_U1-Pad1_ adc_bridge_1		
U4  Net-_U1-Pad2_ pwm dac_bridge_1		
v1  clk GND pulse		
v2  Vin GND DC		
L1  Vin Net-_D1-Pad1_ 100u		
Q1  Net-_D1-Pad1_ pwm GND eSim_NPN		
C1  Vout GND 100u		
R1  Vout GND 100		
U7  Vout plot_v1		
U5  pwm plot_v1		
U2  clk plot_v1		
U6  Vin plot_v1		
D1  Net-_D1-Pad1_ Vout eSim_Diode		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ yt_pwm		

.end
